module d_register (D, clk, Q);
	input D, clk;
	output Q;
	reg Q;
	
	always @(posedge clk)
		Q <= D;
		
endmodule